/*module dff(din, clock, q, qn);
	input din, clock; 
	output reg q, qn; 

	always@(posedge clock)
		begin 
			q = din; 
			qn = ~q; 
		end  
endmodule*/
